Normalizer_2stage.bsv